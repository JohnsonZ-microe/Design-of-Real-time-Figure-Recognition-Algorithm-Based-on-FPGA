library verilog;
use verilog.vl_types.all;
entity gaussian_function_tb is
end gaussian_function_tb;
