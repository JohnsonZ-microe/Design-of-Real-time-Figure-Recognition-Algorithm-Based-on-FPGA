library verilog;
use verilog.vl_types.all;
entity delay_tb is
end delay_tb;
